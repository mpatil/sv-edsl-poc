`ifdef MAIN
module lex;
`endif

//`define LEXDEBUG

`define NLSTATE yyprevious = `YYNEWLINE
`define BEGIN yybgin_ptr = 1 +
`define INITIAL 0
`define YYLERR 0
`define YYSTATE (yyestate_ptr - 1)
`define YYTYPE byte unsigned
`define BUFSIZ 4096 
`ifndef YYLMAX 
`define YYLMAX `BUFSIZ
`endif 

`define lex_output(c) $write(c)
`define unput(c) begin yytchar = (c); if(yytchar == "\n") yylineno--; end
`define yymore() (yymorfg=1)
int yyleng;
int yybgin_ptr = 1;

`define YYISARRAY

typedef byte unsigned Bus[$];
Bus yytext;

int yymorfg;
byte yytchar;
int yyin = -1, yyout = -1;

int yylineno = 1;

function int lex_input();
  yytchar = b.Bgetc();
  if (yytchar == 10) yylineno++;
  if (yytchar == `Beof) return 0;
  lex_input = yytchar;
endfunction

task _yyioinit();
    yyin = 0; yyout = 1;
endtask

typedef struct {
    `YYTYPE verify, advance;
} YYWork;

typedef struct {
  int yystoff_ptr;
  int yyother_ptr;
  int yystops_ptr;
} YYSvf;

/* -*- sv -*- File generated by the BNF Converter (bnfc 2.9.6). */
/* Lexer definition for use with lex */
/* This lex file was machine-generated */
`define YY_BUFFER_LENGTH 4096

string YY_PARSED_STRING;
task YY_BUFFER_APPEND(string s);
  s = {YY_PARSED_STRING, s}; //Do something better here!
endtask
task YY_BUFFER_RESET();
  for(int x = 0; x < `YY_BUFFER_LENGTH; x++)
    YY_PARSED_STRING[x] = 0;
endtask

int yy_mylinenumber = 0;
`define STRING_CAST(x)  string'(x)

`define YYINITIAL 2
`define CHAR 4
`define CHARESC 6
`define CHAREND 8
`define STRING 10
`define ESCAPED 12
`define COMMENT 14
`define YYNEWLINE 10
function int yylex();
	automatic int nstr = 0; //int yyprevious;
  if (yyin == -1) yyin = 0;
  if (yyout == -1) yyout = 1;
  while ((nstr = yylook()) >= 0) begin
    case(nstr)
      0: if(yywrap()) return(0);
      1:      	 return `_SEMI;
      2:      	 return `_LBRACE;
      3:      	 return `_RBRACE;
      4:      	 return `_COMMA;
      5:      	 return `_EQ;
      6:      	 return `_LPAREN;
      7:      	 return `_RPAREN;
      8:      	 return `_DSTAR;
      9:      	 return `_STAR;
      10:      	 return `_SLASH;
      11:      	 return `_PERCENT;
      12:      	 return `_PLUS;
      13:      	 return `_MINUS;
      14:      	 return `_AMP;
      15:      	 return `_CARET;
      16:      	 return `_BAR;
      17:      	 return `_DGT;
      18:      	 return `_DLT;
      19:      	 return `_LT;
      20:      	 return `_LDARROW;
      21:      	 return `_GT;
      22:      	 return `_GTEQ;
      23:      	 return `_DEQ;
      24:      	 return `_BANGEQ;
      25:      	 return `_DAMP;
      26:      	 return `_DBAR;
      27:      	 return `_QUESTION;
      28:      	 return `_COLON;
      29:      	 return `_LBRACK;
      30:      	 return `_RBRACK;
      31:      	 return `_BANG;
      32:      	 return `_TILDE;
      33:      	 return `_DPLUS;
      34:      	 return `_DMINUS;
      35:      	 return `_KW_bin;
      36:      	 return `_KW_break;
      37:      	 return `_KW_ceil;
      38:      	 return `_KW_continue;
      39:      	 return `_KW_defined;
      40:      	 return `_KW_else;
      41:      	 return `_KW_elsif;
      42:      	 return `_KW_fatal;
      43:      	 return `_KW_floor;
      44:      	 return `_KW_for;
      45:      	 return `_KW_forever;
      46:      	 return `_KW_function;
      47:      	 return `_KW_hex;
      48:      	 return `_KW_if;
      49:      	 return `_KW_48;
      50:      	 return `_KW_log2;
      51:      	 return `_KW_print;
      52:      	 return `_KW_procedure;
      53:      	 return `_KW_regrd;
      54:      	 return `_KW_regwr;
      55:      	 return `_KW_return;
      56:      	 return `_KW_sys;
      57:      	 return `_KW_var;
      58:      	 return `_KW_wait;
      59:      	 return `_KW_while;
      60: ++yy_mylinenumber;
      61: `BEGIN `COMMENT;
      62: `BEGIN `YYINITIAL;
      63: /* skip */;
      64: ++yy_mylinenumber;
      65:    	 begin  yylval._string = `STRING_CAST(yytext); return `T_Decimal_Number;  end
      66:    	 begin  yylval._string = `STRING_CAST(yytext); return `T_Real_Number;  end
      67:    	 begin  yylval._string = `STRING_CAST(yytext); return `T_BinaryNumber;  end
      68:    	 begin  yylval._string = `STRING_CAST(yytext); return `T_HexNumber;  end
      69:    	 begin  yylval._string = `STRING_CAST(yytext); return `T_AnyChars;  end
      70:      	 begin  yylval._string = `STRING_CAST(yytext); return `_IDENT_;  end
      71:  ++yy_mylinenumber ;
      72:      	 /* ignore white space. */;
      73:      	 return `_ERROR_;
      -1: ;
      default: $display($psprintf("bad switch yylook %d",nstr));
    endcase
  end
  return(0);
endfunction /* end of yylex */

/*# line 113 "C.l"*/
 /* Initialization code. */
task initialize_lexer(int inp); `BEGIN `YYINITIAL; endtask



int yyvstop[] = {
0,
71, 0, 
73, 0, 
72, 73, 0, 
71, 72, 0, 
31, 73, 0, 
73, 0, 
11, 73, 0, 
14, 73, 0, 
6, 73, 0, 
7, 73, 0, 
9, 73, 0, 
12, 73, 0, 
4, 73, 0, 
13, 73, 0, 
10, 73, 0, 
65, 73, 0, 
65, 73, 0, 
28, 73, 0, 
1, 73, 0, 
19, 73, 0, 
5, 73, 0, 
21, 73, 0, 
27, 73, 0, 
70, 73, 0, 
29, 73, 0, 
30, 73, 0, 
15, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
70, 73, 0, 
2, 73, 0, 
16, 73, 0, 
3, 73, 0, 
32, 73, 0, 
63, 0, 
64, 71, 0, 
63, 0, 
24, 0, 
69, 0, 
25, 0, 
8, 0, 
33, 0, 
34, 0, 
61, 0, 
65, 0, 
18, 0, 
20, 0, 
23, 0, 
22, 0, 
17, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
48, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
26, 0, 
62, 0, 
60, 0, 
66, 0, 
67, 0, 
68, 0, 
35, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
44, 70, 0, 
70, 0, 
47, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
56, 70, 0, 
57, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
37, 70, 0, 
70, 0, 
70, 0, 
40, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
50, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
58, 70, 0, 
70, 0, 
36, 70, 0, 
70, 0, 
70, 0, 
41, 70, 0, 
42, 70, 0, 
43, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
51, 70, 0, 
70, 0, 
53, 70, 0, 
54, 70, 0, 
70, 0, 
59, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
70, 0, 
55, 70, 0, 
70, 0, 
39, 70, 0, 
45, 70, 0, 
70, 0, 
70, 0, 
70, 0, 
38, 70, 0, 
46, 70, 0, 
70, 0, 
70, 0, 
49, 70, 0, 
52, 70, 0, 
 0 };

//# define YYTYPE byte unsigned
YYWork yycrank[] = '{
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 3, 18 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 1, 17 },	
 '{ 3, 19 },	 '{ 3, 20 },	 '{ 0, 0 },	 '{ 3, 19 },	
 '{ 65, 0 },	 '{ 65, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 65, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 3, 21 },	 '{ 3, 22 },	 '{ 0, 0 },	 '{ 24, 67 },	
 '{ 3, 23 },	 '{ 3, 24 },	 '{ 3, 18 },	 '{ 3, 25 },	
 '{ 3, 26 },	 '{ 3, 27 },	 '{ 3, 28 },	 '{ 3, 29 },	
 '{ 3, 30 },	 '{ 16, 63 },	 '{ 3, 31 },	 '{ 3, 32 },	
 '{ 3, 33 },	 '{ 3, 33 },	 '{ 3, 33 },	 '{ 3, 33 },	
 '{ 3, 33 },	 '{ 3, 33 },	 '{ 3, 33 },	 '{ 3, 33 },	
 '{ 3, 33 },	 '{ 3, 34 },	 '{ 3, 35 },	 '{ 3, 36 },	
 '{ 3, 37 },	 '{ 3, 38 },	 '{ 3, 39 },	 '{ 21, 64 },	
 '{ 3, 40 },	 '{ 27, 68 },	 '{ 28, 69 },	 '{ 30, 70 },	
 '{ 31, 71 },	 '{ 36, 77 },	 '{ 36, 78 },	 '{ 37, 79 },	
 '{ 33, 73 },	 '{ 31, 72 },	 '{ 33, 74 },	 '{ 33, 74 },	
 '{ 33, 74 },	 '{ 33, 74 },	 '{ 33, 74 },	 '{ 33, 74 },	
 '{ 33, 74 },	 '{ 33, 74 },	 '{ 33, 74 },	 '{ 33, 74 },	
 '{ 38, 80 },	 '{ 38, 81 },	 '{ 63, 104 },	 '{ 75, 107 },	
 '{ 75, 107 },	 '{ 121, 141 },	 '{ 3, 41 },	 '{ 0, 0 },	
 '{ 3, 42 },	 '{ 3, 43 },	 '{ 55, 100 },	 '{ 107, 107 },	
 '{ 108, 108 },	 '{ 3, 44 },	 '{ 3, 45 },	 '{ 3, 46 },	
 '{ 3, 47 },	 '{ 3, 48 },	 '{ 45, 85 },	 '{ 3, 49 },	
 '{ 3, 50 },	 '{ 46, 87 },	 '{ 44, 83 },	 '{ 3, 51 },	
 '{ 47, 88 },	 '{ 49, 93 },	 '{ 51, 96 },	 '{ 3, 52 },	
 '{ 45, 86 },	 '{ 3, 53 },	 '{ 3, 54 },	 '{ 44, 84 },	
 '{ 52, 97 },	 '{ 3, 55 },	 '{ 3, 56 },	 '{ 50, 94 },	
 '{ 53, 98 },	 '{ 54, 99 },	 '{ 3, 57 },	 '{ 3, 58 },	
 '{ 3, 59 },	 '{ 3, 60 },	 '{ 4, 21 },	 '{ 50, 95 },	
 '{ 58, 103 },	 '{ 83, 109 },	 '{ 4, 23 },	 '{ 4, 24 },	
 '{ 56, 101 },	 '{ 4, 25 },	 '{ 4, 26 },	 '{ 4, 27 },	
 '{ 4, 28 },	 '{ 4, 29 },	 '{ 4, 30 },	 '{ 56, 102 },	
 '{ 4, 31 },	 '{ 84, 110 },	 '{ 4, 33 },	 '{ 4, 33 },	
 '{ 4, 33 },	 '{ 4, 33 },	 '{ 4, 33 },	 '{ 4, 33 },	
 '{ 4, 33 },	 '{ 4, 33 },	 '{ 4, 33 },	 '{ 4, 34 },	
 '{ 4, 35 },	 '{ 4, 36 },	 '{ 4, 37 },	 '{ 4, 38 },	
 '{ 4, 39 },	 '{ 85, 111 },	 '{ 86, 112 },	 '{ 87, 113 },	
 '{ 88, 114 },	 '{ 89, 115 },	 '{ 32, 73 },	 '{ 48, 89 },	
 '{ 32, 74 },	 '{ 32, 74 },	 '{ 32, 74 },	 '{ 32, 74 },	
 '{ 32, 74 },	 '{ 32, 74 },	 '{ 32, 74 },	 '{ 32, 74 },	
 '{ 32, 74 },	 '{ 32, 74 },	 '{ 48, 90 },	 '{ 90, 116 },	
 '{ 91, 117 },	 '{ 48, 91 },	 '{ 92, 118 },	 '{ 93, 119 },	
 '{ 95, 120 },	 '{ 96, 121 },	 '{ 32, 75 },	 '{ 48, 92 },	
 '{ 4, 41 },	 '{ 99, 126 },	 '{ 4, 42 },	 '{ 4, 43 },	
 '{ 100, 127 },	 '{ 98, 124 },	 '{ 97, 122 },	 '{ 4, 44 },	
 '{ 4, 45 },	 '{ 4, 46 },	 '{ 4, 47 },	 '{ 4, 48 },	
 '{ 97, 123 },	 '{ 4, 49 },	 '{ 4, 50 },	 '{ 101, 128 },	
 '{ 102, 129 },	 '{ 4, 51 },	 '{ 98, 125 },	 '{ 110, 130 },	
 '{ 32, 76 },	 '{ 4, 52 },	 '{ 111, 131 },	 '{ 4, 53 },	
 '{ 4, 54 },	 '{ 112, 132 },	 '{ 113, 133 },	 '{ 4, 55 },	
 '{ 4, 56 },	 '{ 15, 61 },	 '{ 32, 75 },	 '{ 115, 136 },	
 '{ 4, 57 },	 '{ 4, 58 },	 '{ 4, 59 },	 '{ 4, 60 },	
 '{ 22, 65 },	 '{ 15, 61 },	 '{ 15, 62 },	 '{ 114, 134 },	
 '{ 15, 61 },	 '{ 116, 137 },	 '{ 117, 138 },	 '{ 114, 135 },	
 '{ 22, 0 },	 '{ 22, 0 },	 '{ 118, 139 },	 '{ 22, 65 },	
 '{ 22, 0 },	 '{ 72, 72 },	 '{ 120, 140 },	 '{ 122, 142 },	
 '{ 32, 76 },	 '{ 123, 143 },	 '{ 124, 144 },	 '{ 125, 146 },	
 '{ 128, 147 },	 '{ 72, 72 },	 '{ 72, 105 },	 '{ 124, 145 },	
 '{ 72, 72 },	 '{ 129, 148 },	 '{ 15, 61 },	 '{ 130, 149 },	
 '{ 132, 150 },	 '{ 133, 151 },	 '{ 135, 152 },	 '{ 15, 61 },	
 '{ 136, 153 },	 '{ 22, 66 },	 '{ 15, 63 },	 '{ 137, 154 },	
 '{ 138, 155 },	 '{ 139, 156 },	 '{ 22, 65 },	 '{ 140, 157 },	
 '{ 15, 61 },	 '{ 142, 158 },	 '{ 143, 159 },	 '{ 144, 160 },	
 '{ 145, 161 },	 '{ 146, 162 },	 '{ 72, 72 },	 '{ 22, 65 },	
 '{ 148, 163 },	 '{ 150, 164 },	 '{ 151, 165 },	 '{ 72, 72 },	
 '{ 155, 166 },	 '{ 156, 167 },	 '{ 157, 168 },	 '{ 159, 169 },	
 '{ 40, 82 },	 '{ 15, 61 },	 '{ 162, 170 },	 '{ 164, 171 },	
 '{ 72, 72 },	 '{ 165, 172 },	 '{ 166, 173 },	 '{ 167, 174 },	
 '{ 22, 65 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 168, 175 },	
 '{ 169, 176 },	 '{ 72, 72 },	 '{ 171, 177 },	 '{ 174, 178 },	
 '{ 175, 179 },	 '{ 176, 180 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 179, 181 },	 '{ 180, 182 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 40, 82 },	 '{ 0, 0 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	 '{ 40, 82 },	
 '{ 73, 106 },	 '{ 73, 106 },	 '{ 73, 106 },	 '{ 73, 106 },	
 '{ 73, 106 },	 '{ 73, 106 },	 '{ 73, 106 },	 '{ 73, 106 },	
 '{ 73, 106 },	 '{ 73, 106 },	 '{ 76, 108 },	 '{ 76, 108 },	
 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	
 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 76, 108 },	
 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	
 '{ 76, 108 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 76, 108 },	
 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	 '{ 76, 108 },	
 '{ 76, 108 },	 '{ 0, 0 },	 '{ 0, 0 },	 '{ 0, 0 },	
 '{0, 0}};

YYSvf yysvec[] = '{
 '{ 0, 0, 0 },
 '{ 1, 0, 0 },
  /* state 0 */ '{ 0, 1, 0 },
  /* state 1 */ '{ -3, 0, 0 },
  /* state 2 */ '{ -97, 3, 0 },
  /* state 3 */ '{ 0, 1, 0 },
  /* state 4 */ '{ 0, 1, 0 },
  /* state 5 */ '{ 0, 1, 0 },
  /* state 6 */ '{ 0, 1, 0 },
  /* state 7 */ '{ 0, 1, 0 },
  /* state 8 */ '{ 0, 1, 0 },
  /* state 9 */ '{ 0, 1, 0 },
  /* state 10 */ '{ 0, 1, 0 },
  /* state 11 */ '{ 0, 1, 0 },
  /* state 12 */ '{ 0, 1, 0 },
  /* state 13 */ '{ -216, 0, 0 },
  /* state 14 */ '{ -7, 15, 0 },
  /* state 15 */ '{ 0, 0, 1 },
  /* state 16 */ '{ 0, 0, 3 },
  /* state 17 */ '{ 0, 0, 5 },
  /* state 18 */ '{ 0, 0, 8 },
  /* state 19 */ '{ 6, 0, 11 },
  /* state 20 */ '{ -223, 0, 14 },
  /* state 21 */ '{ 0, 0, 16 },
  /* state 22 */ '{ 1, 0, 19 },
  /* state 23 */ '{ 0, 0, 22 },
  /* state 24 */ '{ 0, 0, 25 },
  /* state 25 */ '{ 27, 0, 28 },
  /* state 26 */ '{ 27, 0, 31 },
  /* state 27 */ '{ 0, 0, 34 },
  /* state 28 */ '{ 26, 0, 37 },
  /* state 29 */ '{ 30, 0, 40 },
  /* state 30 */ '{ 120, 0, 43 },
  /* state 31 */ '{ 30, 0, 46 },
  /* state 32 */ '{ 0, 0, 49 },
  /* state 33 */ '{ 0, 0, 52 },
  /* state 34 */ '{ 13, 0, 55 },
  /* state 35 */ '{ 14, 0, 58 },
  /* state 36 */ '{ 27, 0, 61 },
  /* state 37 */ '{ 0, 0, 64 },
  /* state 38 */ '{ 241, 0, 67 },
  /* state 39 */ '{ 0, 0, 70 },
  /* state 40 */ '{ 0, 0, 73 },
  /* state 41 */ '{ 0, 0, 76 },
  /* state 42 */ '{ 5, 40, 79 },
  /* state 43 */ '{ 5, 40, 82 },
  /* state 44 */ '{ 8, 40, 85 },
  /* state 45 */ '{ 4, 40, 88 },
  /* state 46 */ '{ 70, 40, 91 },
  /* state 47 */ '{ 12, 40, 94 },
  /* state 48 */ '{ 21, 40, 97 },
  /* state 49 */ '{ 3, 40, 100 },
  /* state 50 */ '{ 6, 40, 103 },
  /* state 51 */ '{ 23, 40, 106 },
  /* state 52 */ '{ 4, 40, 109 },
  /* state 53 */ '{ 1, 40, 112 },
  /* state 54 */ '{ 39, 40, 115 },
  /* state 55 */ '{ 0, 0, 118 },
  /* state 56 */ '{ 8, 0, 121 },
  /* state 57 */ '{ 0, 0, 124 },
  /* state 58 */ '{ 0, 0, 127 },
  /* state 59 */ '{ 0, 0, 130 },
  /* state 60 */ '{ 0, 0, 132 },
  /* state 61 */ '{ 43, 0, 135 },
  /* state 62 */ '{ 0, 0, 137 },
  /* state 63 */ '{ -7, 22, 0 },
  /* state 64 */ '{ 0, 0, 139 },
  /* state 65 */ '{ 0, 0, 141 },
  /* state 66 */ '{ 0, 0, 143 },
  /* state 67 */ '{ 0, 0, 145 },
  /* state 68 */ '{ 0, 0, 147 },
  /* state 69 */ '{ 0, 0, 149 },
  /* state 70 */ '{ -236, 0, 0 },
  /* state 71 */ '{ 316, 0, 0 },
  /* state 72 */ '{ 0, 33, 151 },
  /* state 73 */ '{ 43, 0, 0 },
  /* state 74 */ '{ 326, 0, 0 },
  /* state 75 */ '{ 0, 0, 153 },
  /* state 76 */ '{ 0, 0, 155 },
  /* state 77 */ '{ 0, 0, 157 },
  /* state 78 */ '{ 0, 0, 159 },
  /* state 79 */ '{ 0, 0, 161 },
  /* state 80 */ '{ 0, 40, 163 },
  /* state 81 */ '{ 23, 40, 165 },
  /* state 82 */ '{ 44, 40, 167 },
  /* state 83 */ '{ 56, 40, 169 },
  /* state 84 */ '{ 52, 40, 171 },
  /* state 85 */ '{ 61, 40, 173 },
  /* state 86 */ '{ 49, 40, 175 },
  /* state 87 */ '{ 49, 40, 177 },
  /* state 88 */ '{ 68, 40, 179 },
  /* state 89 */ '{ 66, 40, 181 },
  /* state 90 */ '{ 72, 40, 183 },
  /* state 91 */ '{ 63, 40, 185 },
  /* state 92 */ '{ 0, 40, 187 },
  /* state 93 */ '{ 68, 40, 190 },
  /* state 94 */ '{ 82, 40, 192 },
  /* state 95 */ '{ 89, 40, 194 },
  /* state 96 */ '{ 90, 40, 196 },
  /* state 97 */ '{ 74, 40, 198 },
  /* state 98 */ '{ 78, 40, 200 },
  /* state 99 */ '{ 98, 40, 202 },
  /* state 100 */ '{ 99, 40, 204 },
  /* state 101 */ '{ 0, 0, 206 },
  /* state 102 */ '{ 0, 0, 208 },
  /* state 103 */ '{ 0, 0, 210 },
  /* state 104 */ '{ 0, 73, 212 },
  /* state 105 */ '{ 4, 75, 214 },
  /* state 106 */ '{ 5, 76, 216 },
  /* state 107 */ '{ 0, 40, 218 },
  /* state 108 */ '{ 110, 40, 221 },
  /* state 109 */ '{ 102, 40, 223 },
  /* state 110 */ '{ 97, 40, 225 },
  /* state 111 */ '{ 109, 40, 227 },
  /* state 112 */ '{ 126, 40, 229 },
  /* state 113 */ '{ 122, 40, 231 },
  /* state 114 */ '{ 118, 40, 233 },
  /* state 115 */ '{ 129, 40, 235 },
  /* state 116 */ '{ 135, 40, 238 },
  /* state 117 */ '{ 0, 40, 240 },
  /* state 118 */ '{ 124, 40, 243 },
  /* state 119 */ '{ 43, 40, 245 },
  /* state 120 */ '{ 129, 40, 247 },
  /* state 121 */ '{ 142, 40, 249 },
  /* state 122 */ '{ 128, 40, 251 },
  /* state 123 */ '{ 126, 40, 253 },
  /* state 124 */ '{ 0, 40, 255 },
  /* state 125 */ '{ 0, 40, 258 },
  /* state 126 */ '{ 128, 40, 261 },
  /* state 127 */ '{ 141, 40, 263 },
  /* state 128 */ '{ 144, 40, 265 },
  /* state 129 */ '{ 0, 40, 267 },
  /* state 130 */ '{ 147, 40, 270 },
  /* state 131 */ '{ 143, 40, 272 },
  /* state 132 */ '{ 0, 40, 274 },
  /* state 133 */ '{ 152, 40, 277 },
  /* state 134 */ '{ 148, 40, 279 },
  /* state 135 */ '{ 145, 40, 281 },
  /* state 136 */ '{ 142, 40, 283 },
  /* state 137 */ '{ 145, 40, 285 },
  /* state 138 */ '{ 168, 40, 287 },
  /* state 139 */ '{ 0, 40, 289 },
  /* state 140 */ '{ 149, 40, 292 },
  /* state 141 */ '{ 165, 40, 294 },
  /* state 142 */ '{ 167, 40, 296 },
  /* state 143 */ '{ 154, 40, 298 },
  /* state 144 */ '{ 155, 40, 300 },
  /* state 145 */ '{ 0, 40, 302 },
  /* state 146 */ '{ 171, 40, 305 },
  /* state 147 */ '{ 0, 40, 307 },
  /* state 148 */ '{ 163, 40, 310 },
  /* state 149 */ '{ 173, 40, 312 },
  /* state 150 */ '{ 0, 40, 314 },
  /* state 151 */ '{ 0, 40, 317 },
  /* state 152 */ '{ 0, 40, 320 },
  /* state 153 */ '{ 175, 40, 323 },
  /* state 154 */ '{ 172, 40, 325 },
  /* state 155 */ '{ 159, 40, 327 },
  /* state 156 */ '{ 0, 40, 329 },
  /* state 157 */ '{ 179, 40, 332 },
  /* state 158 */ '{ 0, 40, 334 },
  /* state 159 */ '{ 0, 40, 337 },
  /* state 160 */ '{ 172, 40, 340 },
  /* state 161 */ '{ 0, 40, 342 },
  /* state 162 */ '{ 166, 40, 345 },
  /* state 163 */ '{ 185, 40, 347 },
  /* state 164 */ '{ 172, 40, 349 },
  /* state 165 */ '{ 176, 40, 351 },
  /* state 166 */ '{ 202, 40, 353 },
  /* state 167 */ '{ 183, 40, 355 },
  /* state 168 */ '{ 0, 40, 357 },
  /* state 169 */ '{ 201, 40, 360 },
  /* state 170 */ '{ 0, 40, 362 },
  /* state 171 */ '{ 0, 40, 365 },
  /* state 172 */ '{ 193, 40, 368 },
  /* state 173 */ '{ 199, 40, 370 },
  /* state 174 */ '{ 191, 40, 372 },
  /* state 175 */ '{ 0, 40, 374 },
  /* state 176 */ '{ 0, 40, 377 },
  /* state 177 */ '{ 216, 40, 380 },
  /* state 178 */ '{ 232, 40, 382 },
  /* state 179 */ '{ 0, 40, 384 },
  /* state 180 */ '{ 0, 40, 387 },
  /* state 181 */ '{ 0, 0, 0}
};

int yytop_ptr = 428;
//int yybgin_ptr = 1;
byte unsigned yymatch[] = {
  0,   1,   1,   1,   1,   1,   1,   1, 
  1,   9,  10,   1,  12,   9,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
 12,   1,  34,   1,   1,   1,   1,  39, 
  1,   1,   1,   1,   1,   1,   1,   1, 
 48,  48,  48,  48,  48,  48,  48,  48, 
 48,  48,   1,   1,   1,   1,   1,   1, 
  1,  65,  65,  65,  65,  65,  65,  65, 
 65,  65,  65,  65,  65,  65,  65,  65, 
 65,  65,  65,  65,  65,  65,  65,  65, 
 65,  65,  65,   1,   1,   1,   1,  39, 
  1,  65,  65,  65,  65,  65,  65,  65, 
 65,  65,  65,  65,  65,  65,  65,  65, 
 65,  65,  65,  65,  65,  65,  65,  65, 
 65,  65,  65,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
  1,   1,   1,   1,   1,   1,   1,   1, 
0 };

byte unsigned yyextra[] = {
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,
 0 };

`define NLSTATE yyprevious = `YYNEWLINE

int yylstate[`YYLMAX];

int yylstate_ptr, yylsp_ptr, yyolsp_ptr;

int yyfnd_ptr;
int yyestate_ptr;
int yyprevious = `YYNEWLINE;

task allprint(byte c);
  case(c)
    "\n": $write("\\n");
    "\t": $write("\\t");
    "\b": $write("\\b");
    " " : $write("\\\bb");
    default: $write($psprintf("%s",c));
  endcase
  return;
endtask

task sprint(string pc);
  $write($psprintf("%s", pc));
endtask

function int yylook();
  int yystate_ptr, lsp_ptr;
  int yyt_ptr;
  int yyz_ptr;
  byte unsigned yych;
  int yyfirst;
  int yyr_ptr;

  int debug;

  int yylastch_ptr;

  /* start off machines */
`ifdef LEXDEBUG
  debug = 1;
`endif

  yyfirst = 1;

  if (!yymorfg) begin
    yylastch_ptr = 0;
    //yytext = {};
  end
  else begin
    yymorfg = 0;
    yylastch_ptr = yyleng;
  end

  forever begin
`ifdef LEXDEBUG
    $write ("\n\nouter yylastch_ptr = %0d yyleng = %0d yytext[0] = %0d\n", yylastch_ptr, yyleng, yytext[0]);
`endif
    lsp_ptr = 0;

    yyestate_ptr = yybgin_ptr;
    yystate_ptr = yybgin_ptr;

    if (yyprevious == `YYNEWLINE) yystate_ptr++;

    forever begin
      automatic bit tryagain = 0;
      automatic bit contin = 0;

`ifdef LEXDEBUG
      if (debug) $write ($psprintf("state %0d\n", yystate_ptr - 1));
`endif

      yyt_ptr = yysvec[yystate_ptr].yystoff_ptr;

      if (yyt_ptr == 0 && !yyfirst) begin  /* may not be any transitions */
`ifdef LEXDEBUG
        $write ("\n\nbreaking\n");
`endif
        yyz_ptr = yysvec[yystate_ptr].yyother_ptr;
        if (yyz_ptr == 0) break;
        if (yysvec[yyz_ptr].yystoff_ptr == 0) break;
      end

      yych = lex_input();
      begin
        yytext[yylastch_ptr]  = yych;
`ifdef LEXDEBUG
        $write("yytext: %p\n", yytext);
        $write("yytext: %s\n", string'(yytext));
`endif
      end
      yylastch_ptr++;

`ifdef LEXDEBUG
      $write("len: %0d yych = %0d yytext: %s yylastch_ptr: %0d\n", yytext.size(), yych, string'(yytext), yylastch_ptr);
`endif

      if (yylastch_ptr > `YYLMAX) begin
        $write($psprintf("Input string too long, limit %d\n", `YYLMAX));
        $fatal(1);
      end
      yyfirst = 0;

      do begin : try_again
        contin = 0;
`ifdef LEXDEBUG
        if (debug) begin
          $write("char ");
          allprint(yych);
          $write("\n");
        end
        $write("yyt = %0d yyr = %0d yytop = %0d yytext = %s\n", yyt_ptr, yyr_ptr, yytop_ptr, string'(yytext));
`endif
        yyr_ptr = yyt_ptr;
        if ( yyt_ptr > 0) begin
          yyt_ptr = yyr_ptr + yych;
`ifdef LEXDEBUG
          $write(">yyt = %0d yytop = %0d yystate = %0d\n", yyt_ptr, yytop_ptr, yystate_ptr);
`endif
          if (yyt_ptr <= yytop_ptr && yycrank[yyt_ptr].verify == yystate_ptr) begin
            if (yycrank[yyt_ptr].advance == `YYLERR) begin   /* error transitions */
`ifdef LEXDEBUG
              $write(">unput\n");
`endif
              `unput(yytext[--yylastch_ptr]);
              break;
            end
            yystate_ptr = yycrank[yyt_ptr].advance;
            yylstate[lsp_ptr++] = yystate_ptr;
`ifdef LEXDEBUG
            $write("yystate = %0d\n", yystate_ptr);
`endif
            if (lsp_ptr > `YYLMAX) begin
              $write($psprintf("Input string too long, limit %d\n", `YYLMAX));
              $fatal(1);
            end
`ifdef LEXDEBUG
            if (debug) begin
              $write( $psprintf("+\nstate %0d char ", yystate_ptr - 1));
              allprint(yych);
              $write("\n");
            end
`endif
            contin = 1;
            break;
          end
        end
        else if (yyt_ptr < 0) begin    /* r < yycrank */
          yyr_ptr = -1 * yyt_ptr;
          yyt_ptr = yyr_ptr;
`ifdef LEXDEBUG
          if (debug) $write("compressed state\n");
`endif
          yyt_ptr = yyt_ptr + yych;
`ifdef LEXDEBUG
          $write("yyt = %0d yyr = %0d\n", yyt_ptr, yyr_ptr);
`endif
          if (yyt_ptr <= yytop_ptr && yycrank[yyt_ptr].verify == yystate_ptr) begin
            if (yycrank[yyt_ptr].advance == `YYLERR) begin    /* error transitions */
`ifdef LEXDEBUG
              $write(">>unput\n");
`endif
              `unput(yytext[--yylastch_ptr]);
              break;
            end
            yystate_ptr = yycrank[yyt_ptr].advance;
            yylstate[lsp_ptr++] = yystate_ptr;
            if (lsp_ptr > `YYLMAX) begin
              $write($psprintf("Input string too long, limit %d\n", `YYLMAX));
              $fatal(1);
            end
`ifdef LEXDEBUG
            if (debug) begin
              $write( $psprintf("++\nstate %0d char ", yystate_ptr - 1));
              allprint(yych);
              $write("\n");
            end
`endif
            contin = 1;
            break;
          end
          yyt_ptr = yyr_ptr + yymatch[yych];
`ifdef LEXDEBUG
          if (debug) begin
            $write ("try fall back character ");
            allprint(yymatch[yych]);
            $write("\n");
          end
          $write("yyt = %0d yyr = %0d\n", yyt_ptr, yyr_ptr);
`endif
          if (yyt_ptr <= yytop_ptr && yycrank[yyt_ptr].verify == yystate_ptr) begin
            if (yycrank[yyt_ptr].advance == `YYLERR) begin   /* error transition */
`ifdef LEXDEBUG
              $write(">>>unput\n");
`endif
              `unput(yytext[--yylastch_ptr]);
              break;
            end
            yystate_ptr = yycrank[yyt_ptr].advance;
            yylstate[lsp_ptr++] = yystate_ptr;
            if (lsp_ptr > `YYLMAX) begin
              $write($psprintf("Input string too long, limit %d\n", `YYLMAX));
              $fatal(1);
            end
`ifdef LEXDEBUG
            if (debug) begin
              $write( $psprintf("+++\nstate %0d char ", yystate_ptr - 1));
              allprint(yych);
              $write("\n");
            end
`endif
            contin = 1;
            break;
          end
        end
        yystate_ptr = yysvec[yystate_ptr].yyother_ptr;
        if (yystate_ptr)
          yyt_ptr = yysvec[yystate_ptr].yystoff_ptr;
        tryagain = yystate_ptr && yyt_ptr;

        if (tryagain) begin
`ifdef LEXDEBUG
          if(debug) $write($psprintf("fall back to state %0d\n", yystate_ptr - 1));
          $write("--yyt = %0d yyr = %0d\n", yyt_ptr, yyr_ptr);
`endif
        end
      end while(tryagain);
 
      if (contin) begin
`ifdef LEXDEBUG
        $write("here\n")
`endif
        ;
      end else begin
`ifdef LEXDEBUG
        $write(">>>>unput\n");
`endif
        `unput(yytext[--yylastch_ptr]);
        b.Bungetc();
        break;
      end
    end
`ifdef LEXDEBUG
    if (debug) begin
      $write($psprintf("stopped at %0d with ", yylstate[lsp_ptr - 1] - 1));
      allprint(yych);
      $write("\n");
    end
    $write($psprintf("lsp: %0d\n", lsp_ptr));
`endif
    while (lsp_ptr-- > 0) begin
      yytext[yylastch_ptr--] = 0;
`ifdef LEXDEBUG
      $write($psprintf("lsp: %0d yyfnd: %0d next yyfnd: %0d yytext: %s\n", lsp_ptr, yyfnd_ptr, yysvec[yylstate[lsp_ptr]].yystops_ptr, string'(yytext)));
`endif
      if (yylstate[lsp_ptr] != 0)
        yyfnd_ptr = yysvec[yylstate[lsp_ptr]].yystops_ptr;
      if (yyfnd_ptr > 0) begin
        yyolsp_ptr = lsp_ptr;
`ifdef LEXDEBUG
        $write($psprintf("yyextra[%0d] = %0d\n", yyvstop[yyfnd_ptr], yyextra[yyvstop[yyfnd_ptr]]));
`endif
        if (yyextra[yyvstop[yyfnd_ptr]]) begin        /* must backup */
          while(yyback(yysvec[yylstate[lsp_ptr]].yystops_ptr, -1 * yyfnd_ptr) != 1 && lsp_ptr > 0)begin
            lsp_ptr--;
`ifdef LEXDEBUG
            $write(">>>>>unput\n");
`endif
            `unput(yytext[yylastch_ptr--]);
          end
        end
        yyprevious = yytext[yylastch_ptr];
        yylsp_ptr = lsp_ptr;
        yyleng = yylastch_ptr + 1;
        yytext = yytext[0:yyleng - 1];
`ifdef LEXDEBUG
        if(debug) begin
          $write("\nmatch ");
          $write(" (yyleng: %0d, yylastch_ptr: %0d) ", yyleng, yylastch_ptr);
          $write("%s", string'(yytext));
          $write($psprintf(" action %0d\n\n", yyvstop[yyfnd_ptr]));
        end
`endif
        return(yyvstop[yyfnd_ptr++]); // XXX
      end
`ifdef LEXDEBUG
      $write(">>>>>>unput\n");
`endif
      `unput(yytext[yylastch_ptr]);
    end
    if (yytext[0] == 0  /* && feof(yyin) */)
    begin
      if(debug) $write("Exiting\n");
      return(0);
    end
    yyprevious = lex_input();
    yytext[0] = yyprevious;
    if (yyprevious > 0)
      `lex_output(yyprevious);
    yytext = {};
    yylastch_ptr = 0;
`ifdef LEXDEBUG
    if(debug) $write("\n");
`endif
  end
endfunction

function int yyback(int p, int m);
  if (yyvstop[p]==0) return(0);
  while (yyvstop[p]) begin
    if (yyvstop[p++] == m)
      return(1);
  end
  return(0);
endfunction

/* the following are only used in the lex library */
function int yyinput();
  return(lex_input());
endfunction

task  yyoutput(int c);
  `lex_output(c);
endtask

task yyunput(int c);
  `unput(c);
endtask

`ifdef MAIN
initial begin
  string filename;
  int tok;

  if ($value$plusargs("input=%s", filename))
    b = Bopen(filename, `OREAD);

  $write("\n");
  initialize_lexer(0);
  tok = yylex();
  while(tok) begin
    $write($psprintf("token: %0d\n", tok));
    tok = yylex();
  end
  $write($psprintf("token: %0d\n", tok));
  $write("\n");
end
endmodule
`endif
